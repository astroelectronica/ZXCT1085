.title KiCad schematic
.include "C:/AE/ZXCT1085/_models/C2012CH2W101J060AA_p.mod"
.include "C:/AE/ZXCT1085/_models/C2012X7R2A104K125AA_p.mod"
.include "C:/AE/ZXCT1085/_models/ZXCT1085E5TA.LIB"
XU2 VDD 0 C2012X7R2A104K125AA_p
R5 /VOCM 0 {RPD}
XU1 /VOCM 0 /VIN /SN VDD ZXCT1085E5TA
V2 VDD 0 DC {VSUPPLY} 
R2 /VIN /VOUT {RSNS}
R1 /VIN /VOUT {RSNS}
V1 /VIN 0 DC {VSOURCE} 
R3 /VOUT /SN {RN}
XU3 /VIN /SN C2012CH2W101J060AA_p
I1 /VOUT 0 DC {ILOAD} 
.end
